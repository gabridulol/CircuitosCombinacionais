`include "./Verilog/Codificador.v"

module Display (
    ports
);
    
endmodule